module State_machine();

endmodule

